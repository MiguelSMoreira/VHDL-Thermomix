----------------------------------------------------------------------------------
-- Company: IST
-- Engineer: Miguel Moreira e Pedro Coimbra
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
--Ficheiro rom_memory_tabela.vhd

--Declaracao das Bibliotecas
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--Declaracao da Entidade
entity rom_memory_tabela is
    Port ( 
            address : in  STD_LOGIC_VECTOR (7 downto 0);
            data : out  STD_LOGIC_VECTOR (44 downto 0)
         );
end rom_memory_tabela;

--Declaracao da arquitectura do Componente
architecture Behavioral of rom_memory_tabela is

  type ram_type is array (0 to 127) 
	 of std_logic_vector(44 downto 0);
	 
	 constant InitValue: ram_type := (
      0 => "00000001" & "00000011" & "000001000000" & "00100000" & "00000010" & "1", --(do bit mais significativo (esquerda) para o bit menos significativo (direita))
		1 => "00000001" & "00000010" & "000000100000" & "00000101" & "00010010" & "0",
		2 => "00000001" & "00000001" & "000000010101" & "00000101" & "00000111" & "1",
		3 => "00000001" & "00000000" & "000000010000" & "00010000" & "00001000" & "0",
		4 => "00000010" & "00000001" & "000000010000" & "00000101" & "00000101" & "1",
		5 => "00000010" & "00000000" & "000000000101" & "00000101" & "00010000" & "0",
		6 => "00000011" & "00000010" & "000001100000" & "00110000" & "00001000" & "1",
		7 => "00000011" & "00000001" & "000000110000" & "00010000" & "00010011" & "1",
		8 => "00000011" & "00000000" & "000000100000" & "00100000" & "00000101" & "0",
		9 => "00000100" & "00000000" & "000010011001" & "10011001" & "00010000" & "0",
		10 => "00000101" & "00001000" & "001001100000" & "01010000" & "00000111" & "0",
		11 => "00000101" & "00000111" & "001000010000" & "00110000" & "00001000" & "1",
		12 => "00000101" & "00000110" & "000110000000" & "01000000" & "00001001" & "0",
		13 => "00000101" & "00000101" & "000101100101" & "00010101" & "00010000" & "1",
		14 => "00000101" & "00000100" & "000101000101" & "00100000" & "00000011" & "0",
		15 => "00000101" & "00000011" & "000100100000" & "00100101" & "00000101" & "1",
		16 => "00000101" & "00000010" & "000010010000" & "00110000" & "00000111" & "0",
		17 => "00000101" & "00000001" & "000001010000" & "01000000" & "00000011" & "0",
		18 => "00000101" & "00000000" & "000000010000" & "00010000" & "00000010" & "0",
		19 => "00000110" & "00000001" & "000001010101" & "00110101" & "00000111" & "0",
		20 => "00000110" & "00000000" & "000000100000" & "00100000" & "00000101" & "0",
		21 => "00000111" & "00000000" & "000000010101" & "00010101" & "00010101" & "0",
		22 => "00001000" & "00000010" & "000001100101" & "00010000" & "00010000" & "1",
		23 => "00001000" & "00000001" & "000001010101" & "01000000" & "00000111" & "0",
		24 => "00001000" & "00000000" & "000000010101" & "00010101" & "00000101" & "0",
		25 => "00001001" & "00000011" & "000001100000" & "00110000" & "00000011" & "1",
		26 => "00001001" & "00000010" & "000000110000" & "00010000" & "00010011" & "0",
		27 => "00001001" & "00000001" & "000000100000" & "00000101" & "00000110" & "1",
		28 => "00001001" & "00000000" & "000000010101" & "00010101" & "00001000" & "0",
	others => "000000000000000000000000000000000000000000000" -- (todas os outros enderecos nao indicados anteriormente)
	);       
 
signal Content_d_mem: ram_type:= InitValue;

begin

data <= Content_d_mem(CONV_INTEGER(address));

end Behavioral;